module mux4to1ifelse(w,s,out);
           input [0:3] w;
           input [1:0] s; // here 1 is MSB and 0 is lsb, so if you write [0:1] , then 
           // for s == 1, it would consider s[0] as MSB and s[1] as LSB. So s = = 1 decimal
           // will be got when s[0] = 0 and s[1] = 1. be careful about this point
           // w can be written both as [3:0] or [0:3] because there is no need for binary to decimal 
           // conversion, thus no need for the concept of MSB or LSB, it is directly assigned 
           // in the always block
           output reg out;
           always @(s) // omitted the dependency on the input
           begin
                     out = w[3]; // omitted one extra else line
                     if(s == 0)
                        out = w[0];
                     else if (s == 1)
                        out = w[1];
                     else if (s == 2)
                        out = w[2];
           end
endmodule