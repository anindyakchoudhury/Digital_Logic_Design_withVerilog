module ternarysystem